--AXI tb from https://github.com/frobino/axi_custom_ip_tb/blob/master/led_controller_1.0/hdl/testbench.vhd

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
library UNISIM;
use UNISIM.VCOMPONENTS.ALL;
entity tb is
 
end tb;

architecture STRUCTURE of tb is

	component xgbe is 
	generic (
		C_S_AXI_DATA_WIDTH	: integer	:= 32;
		C_S_AXI_ADDR_WIDTH	: integer	:= 4
	);
	port (
		clk_156_25MHz	: in std_logic;
		rst_clk_156_25MHz : in std_logic;
		clk_20MHz	: in std_logic;
		rst_clk_20MHz	: in std_logic;

		interrupt	: out std_logic;

		s_axi_aclk	: in std_logic;
		s_axi_aresetn	: in std_logic;
		s_axi_awaddr	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		s_axi_awprot	: in std_logic_vector(2 downto 0);
		s_axi_awvalid	: in std_logic;
		s_axi_awready	: out std_logic;
		s_axi_wdata	: in std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		s_axi_wstrb	: in std_logic_vector((C_S_AXI_DATA_WIDTH/8)-1 downto 0);
		s_axi_wvalid	: in std_logic;
		s_axi_wready	: out std_logic;
		s_axi_bresp	: out std_logic_vector(1 downto 0);
		s_axi_bvalid	: out std_logic;
		s_axi_bready	: in std_logic;
		s_axi_araddr	: in std_logic_vector(C_S_AXI_ADDR_WIDTH-1 downto 0);
		s_axi_arprot	: in std_logic_vector(2 downto 0);
		s_axi_arvalid	: in std_logic;
		s_axi_arready	: out std_logic;
		s_axi_rdata	: out std_logic_vector(C_S_AXI_DATA_WIDTH-1 downto 0);
		s_axi_rresp	: out std_logic_vector(1 downto 0);
		s_axi_rvalid	: out std_logic;
		s_axi_rready	: in std_logic;
		xgmii_rxc : in STD_LOGIC_VECTOR (7 downto 0);
		xgmii_rxd : in STD_LOGIC_VECTOR (63 downto 0);
		xgmii_txc : out STD_LOGIC_VECTOR (7 downto 0);
		xgmii_txd : out STD_LOGIC_VECTOR (63 downto 0);
		xgmii_tx_clk : in std_logic;
		xgmii_rx_clk : in std_logic		
	);
end component xgbe;

  signal xgmii_tx_clk, xgmii_rx_clk : std_logic := '0';
  signal clk_156_25MHz, clk_20MHz, rst_clk_156_25MHz, rst_clk_20MHz : std_logic := '0';
  signal interrupt : std_logic := '0';
  signal s_axi_aclk, s_axi_aresetn, s_axi_arready, s_axi_arvalid, s_axi_awready, s_axi_awvalid : std_logic := '0';
  signal s_axi_bready, s_axi_bvalid, s_axi_rready, s_axi_rvalid, s_axi_wready, s_axi_wvalid : std_logic := '0';
  signal s_axi_rdata, s_axi_wdata : std_logic_vector(31 downto 0) := (others => '0');
  signal s_axi_araddr, s_axi_awaddr, s_axi_wstrb : std_logic_vector(3 downto 0) := (others => '0');
  signal s_axi_arprot, s_axi_awprot : std_logic_vector(2 downto 0) := (others => '0');
  signal s_axi_bresp, s_axi_rresp : std_logic_vector(1 downto 0) := (others => '0');
  
  signal xgmii_rxd, xgmii_txd : std_logic_vector(63 downto 0) := (others => '0');
  signal xgmii_rxc, xgmii_txc : std_logic_vector(7 downto 0) := (others => '0');

  signal ReadIt, SendIt : std_logic := '0';
begin

block_design_i: xgbe
     port map (
	clk_156_25MHz => clk_156_25MHz,
	rst_clk_156_25MHz => rst_clk_156_25MHz,
	clk_20MHz => clk_20MHz,
	rst_clk_20MHz => rst_clk_20MHz,

      interrupt => interrupt,

      s_axi_aclk => s_axi_aclk,
      s_axi_araddr(3 downto 0) => s_axi_araddr(3 downto 0),
      s_axi_aresetn => s_axi_aresetn,
      s_axi_arprot(2 downto 0) => s_axi_arprot(2 downto 0),
      s_axi_arready => s_axi_arready,
      s_axi_arvalid => s_axi_arvalid,
      s_axi_awaddr(3 downto 0) => s_axi_awaddr(3 downto 0),
      s_axi_awprot(2 downto 0) => s_axi_awprot(2 downto 0),
      s_axi_awready => s_axi_awready,
      s_axi_awvalid => s_axi_awvalid,
      s_axi_bready => s_axi_bready,
      s_axi_bresp(1 downto 0) => s_axi_bresp(1 downto 0),
      s_axi_bvalid => s_axi_bvalid,
      s_axi_rdata(31 downto 0) => s_axi_rdata(31 downto 0),
      s_axi_rready => s_axi_rready,
      s_axi_rresp(1 downto 0) => s_axi_rresp(1 downto 0),
      s_axi_rvalid => s_axi_rvalid,
      s_axi_wdata(31 downto 0) => s_axi_wdata(31 downto 0),
      s_axi_wready => s_axi_wready,
      s_axi_wstrb(3 downto 0) => s_axi_wstrb(3 downto 0),
      s_axi_wvalid => s_axi_wvalid,
      xgmii_rxd => xgmii_rxd,
      xgmii_txd => xgmii_txd,
      xgmii_rxc => xgmii_rxc,
      xgmii_txc => xgmii_txc,
      xgmii_tx_clk => xgmii_tx_clk,
      xgmii_rx_clk => xgmii_rx_clk
);

process begin
	wait for 1 ns;
	while true loop
		xgmii_tx_clk <= '0';
		wait for 3.2 ns;
		xgmii_tx_clk <= '1';
		wait for 3.2 ns;
	end loop;
end process;

process begin
	wait for 1.3 ns;
	while true loop
		xgmii_rx_clk <= '1';
		wait for 3.2 ns;
		xgmii_rx_clk <= '0';
		wait for 3.2 ns;
	end loop;
end process;

process begin
    s_axi_aclk <= '0';
    wait for 5 ns;
    s_axi_aclk <= '1';
    wait for 5 ns;
end process;
 
process begin
	clk_156_25MHz <= '1';
	wait for 3.2 ns;
	clk_156_25MHz <= '0';
	wait for 3.2 ns;
end process;

process begin
	clk_20MHz <= '1';
	wait for 25 ns;
	clk_20MHz <= '0';
	wait for 25 ns;
end process;

process begin
	s_axi_aresetn <= '0';
	rst_clk_156_25MHz <= '0';
	rst_clk_20MHz <= '0';
	wait for 6.4 ns;
	rst_clk_156_25MHz <= '1';
	wait for 3.6 ns;
	s_axi_aresetn <= '1';
	wait for 40 ns;
	rst_clk_20MHz <= '1';
	wait;
end process;

send : process
 begin
    s_axi_awvalid<='0';
    s_axi_wvalid<='0';
    s_axi_bready<='0';
    loop
        wait until sendit = '1';
        wait until s_axi_aclk= '0';
            s_axi_awvalid<='1';
            s_axi_wvalid<='1';
        wait until (s_axi_awready and s_axi_wready) = '1';  --client ready to read address/data        
            s_axi_bready<='1';
        wait until s_axi_bvalid = '1';  -- write result valid
            assert s_axi_bresp = "00" report "axi data not written" severity failure;
            s_axi_awvalid<='0';
            s_axi_wvalid<='0';
            s_axi_bready<='1';
        wait until s_axi_bvalid = '0';  -- all finished
            s_axi_bready<='0';
    end loop;
 end process send;

 read : process
  begin
    s_axi_arvalid<='0';
    s_axi_rready<='0';
     loop
         wait until readit = '1';
         wait until s_axi_aclk= '0';
             s_axi_arvalid<='1';
            wait until (s_axi_rvalid) = '1';  --client provided data (removed and s_axi_arready???)
            s_axi_rready<='1';
            s_axi_arvalid <= '0';
            assert s_axi_rresp = "00" report "axi data not written" severity failure;
            wait until (s_axi_rvalid) = '0';
            s_axi_rready<='0';
     end loop;
  end process read;
      
tb : process
begin

	wait until rst_clk_20MHz = '1';

for j in 0 to 1500 loop
	xgmii_rxd <= x"0707070707070707";
	xgmii_rxc <= x"ff";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"d5555555555555fb";
	xgmii_rxc <= x"01";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"0001001000000100";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"88b5000194000002";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000000ffffff00";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000001ffffff01";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000002ffffff02";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000003ffffff03";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000004ffffff04";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"f0000005ffffff05";
	xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
    xgmii_rxd <= x"f0000006ffffff06";
    xgmii_rxc <= x"00";
    wait until rising_edge(clk_156_25MHz);
    xgmii_rxd <= x"f0000007ffffff07";
    xgmii_rxc <= x"00";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"0707fd79d45b7708";
	xgmii_rxc <= x"e0";
	wait until rising_edge(clk_156_25MHz);
	xgmii_rxd <= x"0707070707070707";
	xgmii_rxc <= x"ff";
	wait until rising_edge(clk_156_25MHz);
	end loop;
    
    s_axi_awaddr<="1000";
    s_axi_wdata<=x"00000001";
    s_axi_wstrb<=b"1111";
    sendit<='1';                --start axi write to slave
    wait for 1 ns; 
    sendit<='0'; --clear start send flag
    wait until s_axi_bvalid = '1';
    wait until s_axi_bvalid = '0';  --axi write finished
    s_axi_wstrb<=b"0000";
    
    wait until interrupt = '1';

    s_axi_araddr<="0000";
        readit<='1';                --start axi read from slave
        wait for 1 ns; 
       readit<='0';                --clear "start read" flag
    wait until s_axi_rready = '1';
    wait until s_axi_rready = '0';    --axi_data should be equal to 17
    
    for i in 0 to 50 loop
        s_axi_araddr<="0100";    
        readit<='1';                --start axi read from slave
        wait for 1 ns; 
       readit<='0';                --clear "start read" flag
    wait until s_axi_rready = '1';    --axi_data should be equal to 10000000...
    wait until s_axi_rready = '0';
    end loop; 
    
     
 xgmii_rxd <= x"0707070707070707";
 xgmii_rxc <= x"ff";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"d5555555555555fb";
 xgmii_rxc <= x"01";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"0001001000000100";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"88b5000194000002";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000000ffffff00";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000001ffffff01";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000002ffffff02";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000003ffffff03";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000004ffffff04";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000005ffffff05";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000006ffffff06";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"f0000007ffffff07";
 xgmii_rxc <= x"00";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"0707fd79d45b7708";
 xgmii_rxc <= x"e0";
 wait until rising_edge(clk_156_25MHz);
 xgmii_rxd <= x"0707070707070707";
 xgmii_rxc <= x"ff";
 wait until rising_edge(clk_156_25MHz);
 
  for i in 0 to 50 loop
  s_axi_araddr<="0100";    
  readit<='1';                --start axi read from slave
  wait for 1 ns; 
  readit<='0';                --clear "start read" flag
  wait until s_axi_rready = '1';    --axi_data should be equal to 10000000...
  wait until s_axi_rready = '0';
  end loop; 
    
end process tb;   
     
end structure;
