signal RX_ADDR_STRB, RX_SIZE_STRB, RX_PRCSSD_STRB, RX_PRCSSD_INT 			: std_logic := '0';
signal XGBE_PACKET_RCV	: std_logic := '0';


		RX_ADDR => RX_ADDR,
		RX_ADDR_STRB => RX_ADDR_STRB,
		RX_SIZE => RX_SIZE,
		RX_SIZE_STRB => RX_SIZE_STRB,
		RX_PRCSSD => RX_PRCSSD,
		RX_PRCSSD_STRB => RX_PRCSSD_STRB,
		RX_PRCSSD_INT => RX_PRCSSD_INT,

		XGBE_PACKET_RCV => XGBE_PACKET_RCV,
